//`include "mux.v"

module bs(input [15:0]a, input[3:0]s,input l,output [15:0]b);

wire [15:0]c1,c2,c3;

// l decided the whether arithmetic or logic shift


mux m15(l,a[15],s[0],c1[15]);
mux m14(a[15],a[14],s[0],c1[14]);
mux m13(a[14],a[13],s[0],c1[13]);
mux m12(a[13],a[12],s[0],c1[12]);
mux m11(a[12],a[11],s[0],c1[11]);
mux m10(a[11],a[10],s[0],c1[10]);
mux m9(a[10],a[9],s[0],c1[9]);
mux m8(a[9],a[8],s[0],c1[8]);
mux m7(a[8],a[7],s[0],c1[7]);
mux m6(a[7],a[6],s[0],c1[6]);
mux m5(a[6],a[5],s[0],c1[5]);
mux m4(a[5],a[4],s[0],c1[4]);
mux m3(a[4],a[3],s[0],c1[3]);
mux m2(a[3],a[2],s[0],c1[2]);
mux m1(a[2],a[1],s[0],c1[1]);
mux m0(a[1],a[0],s[0],c1[0]);

mux n15(l,c1[15],s[1],c2[15]);
mux n14(l,c1[14],s[1],c2[14]);
mux n13(c1[15],c1[13],s[1],c2[13]);
mux n12(c1[14],c1[12],s[1],c2[12]);
mux n11(c1[13],c1[11],s[1],c2[11]);
mux n10(c1[12],c1[10],s[1],c2[10]);
mux n9(c1[11],c1[9],s[1],c2[9]);
mux n8(c1[10],c1[8],s[1],c2[8]);
mux n7(c1[9],c1[7],s[1],c2[7]);
mux n6(c1[8],c1[6],s[1],c2[6]);
mux n5(c1[7],c1[5],s[1],c2[5]);
mux n4(c1[6],c1[4],s[1],c2[4]);
mux n3(c1[5],c1[3],s[1],c2[3]);
mux n2(c1[4],c1[2],s[1],c2[2]);
mux n1(c1[3],c1[1],s[1],c2[1]);
mux n0(c1[2],c1[0],s[1],c2[0]);

mux l15(l,c2[15],s[2],c3[15]);
mux l14(l,c2[14],s[2],c3[14]);
mux l13(l,c2[13],s[2],c3[13]);
mux l12(l,c2[12],s[2],c3[12]);
mux l11(c2[15],c2[11],s[2],c3[11]);
mux l10(c2[14],c2[10],s[2],c3[10]);
mux l9(c2[13],c2[9],s[2],c3[9]);
mux l8(c2[12],c2[8],s[2],c3[8]);
mux l7(c2[11],c2[7],s[2],c3[7]);
mux l6(c2[10],c2[6],s[2],c3[6]);
mux l5(c2[9],c2[5],s[2],c3[5]);
mux l4(c2[8],c2[4],s[2],c3[4]);
mux l3(c2[7],c2[3],s[2],c3[3]);
mux l2(c2[6],c2[2],s[2],c3[2]);
mux l1(c2[5],c2[1],s[2],c3[1]);
mux l0(c2[4],c2[0],s[2],c3[0]);

mux o15(l,c3[15],s[3],b[15]);
mux o14(l,c3[14],s[3],b[14]);
mux o13(l,c3[13],s[3],b[13]);
mux o12(l,c3[12],s[3],b[12]);
mux o11(l,c3[11],s[3],b[11]);
mux o10(l,c3[10],s[3],b[10]);
mux o9(l,c3[9],s[3],b[9]);
mux o8(l,c3[8],s[3],b[8]);
mux o7(l,c3[7],s[3],b[7]);
mux o6(c3[15],c3[6],s[3],b[6]);
mux o5(c3[14],c3[5],s[3],b[5]);
mux o4(c3[13],c3[4],s[3],b[4]);
mux o3(c3[12],c3[3],s[3],b[3]);
mux o2(c3[11],c3[2],s[3],b[2]);
mux o1(c3[10],c3[1],s[3],b[1]);
mux o0(c3[9],c3[0],s[3],b[0]);

endmodule 


